LIBRARY ieee;
USE ieee.std_logic_1164.all;

Entity ADDER is
Port( A, B : in std_logic_vector(3 downto 0);
		Ci : in std_logic;
		Co : out std_logic;
		S : out std_logic_vector(3 downto 0));
End ADDER;

ARCHITECTURE structural of ADDER is
Component FA is
Port( A, B, Ci : in std_logic;
		Co, S : out std_logic);
End component;

signal carry : std_logic_vector(3 downto 0);

Begin

U1: FA port map (A => A(0), B=> B(0), Ci => Ci, S => S(0), Co => carry(0));

U2: FA port map (A => A(1), B=> B(1), Ci => carry(0), S => S(1), Co => carry(1));

U3: FA port map (A => A(2), B=> B(2), Ci => carry(1), S => S(2), Co => carry(2));

U4: FA port map (A => A(3), B=> B(3), Ci => carry(2), S => S(3), Co => carry(3));

Co <= carry(3);

End structural;